module NormalCLK (
    outCLK,RST,CLK
);
		input CLK,RST;
		output outCLK;
    //we need 21 DRFF to make clk 5MHZ to 2 HZ
    wire W1,nW1,W2,nW2,W3,nW3,W4,nW4,W5,nW5,W6,nW6,W7,nW7,W8,nW8,W9,nW9,W10,nW10,W11,nW11,W12,nW12,W13,nW13
    ,W14,nW14,W15,nW15,W16,nW16,W17,nW17,W18,nW18,W19,nW19,W20,nW20,nW21;
    DRFF D1(W1,nW1,nW1,RST,CLK);
    DRFF D2(W2,nW2,nW2,RST,W1);
    DRFF D3(W3,nW3,nW3,RST,W2);
    DRFF D4(W4,nW4,nW4,RST,W3);
    DRFF D5(W5,nW5,nW5,RST,W4);
    DRFF D6(W6,nW6,nW6,RST,W5);
    DRFF D7(W7,nW7,nW7,RST,W6);
    DRFF D8(W8,nW8,nW8,RST,W7);
    DRFF D9(W9,nW9,nW9,RST,W8);
    DRFF D10(W10,nW10,nW10,RST,W9);
    DRFF D11(W11,nW11,nW11,RST,W10);
    DRFF D12(W12,nW12,nW12,RST,W11);
    DRFF D13(W13,nW13,nW13,RST,W12);
    DRFF D14(W14,nW14,nW14,RST,W13);
    DRFF D15(W15,nW15,nW15,RST,W14);
    DRFF D16(W16,nW16,nW16,RST,W15);
    DRFF D17(W17,nW17,nW17,RST,W16);
    DRFF D18(W18,nW18,nW18,RST,W17);
    DRFF D19(W19,nW19,nW19,RST,W18);
    DRFF D20(W20,nW20,nW20,RST,W19);
    DRFF D21(outCLK,nW21,nW21,RST,W20);
endmodule